module ratateSignal(
 input clk,
 input [143:0] afterRotate,
 input [143:0] background,
 output canRotate
);

	

endmodule
