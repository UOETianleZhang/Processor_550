module initializer(
	input clk,
	input refresh,
	output [144:0] newShape
);

//parameter [144:0] box = 145'b00001111000000000010;
//parameter [144:0] IShape = 145'd;
parameter [144:0] tShape = 145'h20070;
//parameter [144:0] lShape = 145'd;
//parameter [144:0] zShape = 145'd;

endmodule
